// Options
// `define ERROR_FLAGS 1
`define TWO_STOP_BITS 1
